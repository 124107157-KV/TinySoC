* NGSPICE file created from tiny_soc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

.subckt tiny_soc VGND VPWR clk gpio[0] gpio[1] gpio[2] gpio[3] rst_n uart_rx uart_tx
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_294_ cpu_acc\[4\] _133_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_363_ clknet_3_0__leaf_clk u_cpu.pc_next\[4\] net11 VGND VGND VPWR VPWR cpu_pc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_346_ _056_ _093_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or2_1
X_415_ clknet_3_3__leaf_clk _047_ net14 VGND VGND VPWR VPWR u_cpu.state\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_277_ _055_ _064_ cpu_acc\[2\] VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__o21a_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_200_ net58 _067_ _070_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__o21ai_1
X_329_ net22 _160_ _167_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21o_1
XFILLER_17_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 u_uart.u_tx.bit_cnt\[1\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 u_uart.u_tx.clk_cnt\[0\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ cpu_acc\[4\] _133_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_362_ clknet_3_1__leaf_clk u_cpu.pc_next\[3\] net11 VGND VGND VPWR VPWR cpu_pc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_414_ clknet_3_4__leaf_clk net39 net15 VGND VGND VPWR VPWR u_uart.tx_data\[7\] sky130_fd_sc_hd__dfrtp_1
X_345_ u_uart.tx_start _057_ _083_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ _123_ _125_ cpu_acc\[1\] _116_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ u_uart.tx_data\[5\] net9 net8 u_uart.u_tx.shifter\[6\] VGND VGND VPWR VPWR
+ _167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_259_ net19 _112_ _083_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_5_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout8 _159_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_15_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold20 cpu_acc\[7\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 u_uart.u_tx.clk_cnt\[14\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 cpu_pc\[3\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ cpu_acc\[4\] _133_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ clknet_3_1__leaf_clk u_cpu.pc_next\[2\] net11 VGND VGND VPWR VPWR cpu_pc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_413_ clknet_3_5__leaf_clk _045_ net18 VGND VGND VPWR VPWR u_uart.tx_data\[6\] sky130_fd_sc_hd__dfrtp_1
X_344_ net9 _050_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2b_1
X_275_ _064_ _073_ _116_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__nor3_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_327_ net28 _160_ _166_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a21o_1
X_189_ cpu_acc\[4\] cpu_acc\[5\] cpu_acc\[6\] cpu_acc\[7\] VGND VGND VPWR VPWR _066_
+ sky130_fd_sc_hd__or4_1
X_258_ net10 _111_ _112_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_8_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout9 _158_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
Xhold10 u_uart.u_tx.shifter\[4\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold21 _046_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 u_uart.u_tx.clk_cnt\[6\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 u_uart.u_tx.clk_cnt\[1\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ _124_ _138_ _139_ _116_ net57 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_15_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_360_ clknet_3_1__leaf_clk u_cpu.pc_next\[1\] net14 VGND VGND VPWR VPWR cpu_pc\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ clknet_3_5__leaf_clk _044_ net18 VGND VGND VPWR VPWR u_uart.tx_data\[5\] sky130_fd_sc_hd__dfrtp_1
X_343_ _114_ _115_ _049_ _057_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a31o_1
X_274_ _120_ _121_ _122_ _073_ _065_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__a311o_1
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_326_ u_uart.tx_data\[4\] net9 net8 net22 VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_24_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ u_cpu.state\[1\] _064_ u_cpu.state\[0\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__or3b_1
X_257_ u_uart.u_tx.clk_cnt\[13\] u_uart.u_tx.clk_cnt\[14\] _108_ VGND VGND VPWR VPWR
+ _112_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ cpu_acc\[6\] _116_ _124_ _154_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a22o_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 _029_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 u_uart.tx_data\[4\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 u_uart.u_tx.state\[1\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 cpu_pc\[4\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_290_ _132_ _137_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__or2_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_411_ clknet_3_5__leaf_clk _043_ net18 VGND VGND VPWR VPWR u_uart.tx_data\[4\] sky130_fd_sc_hd__dfrtp_1
X_342_ u_uart.u_tx.state\[0\] _093_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
X_273_ _065_ _073_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__nor2_1
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_325_ net34 _160_ _165_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_256_ u_uart.u_tx.clk_cnt\[13\] _108_ net60 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ _059_ _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_9_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
X_308_ _150_ _153_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__xnor2_1
X_239_ u_uart.u_tx.clk_cnt\[7\] _098_ _100_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__o21a_1
Xhold45 u_uart.u_tx.shifter\[3\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 u_uart.tx_data\[6\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 u_cpu.state\[1\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 u_uart.u_tx.clk_cnt\[12\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_26_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_410_ clknet_3_5__leaf_clk _042_ net15 VGND VGND VPWR VPWR u_uart.tx_data\[3\] sky130_fd_sc_hd__dfrtp_1
X_341_ net9 _171_ _174_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ _120_ _121_ cpu_acc\[0\] VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_324_ u_uart.tx_data\[3\] net9 net8 u_uart.u_tx.shifter\[4\] VGND VGND VPWR VPWR
+ _165_ sky130_fd_sc_hd__a22o_1
X_255_ net56 _108_ _110_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ cpu_pc\[2\] cpu_pc\[3\] VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__or2_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_4
X_307_ _151_ _152_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and2b_1
X_238_ u_uart.u_tx.clk_cnt\[7\] _098_ net10 VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 _048_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 cpu_pc\[5\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 u_uart.u_tx.clk_cnt\[9\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _093_ _115_ _172_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__or3_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_271_ cpu_acc\[0\] _059_ _063_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__or3_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_323_ net21 _160_ _164_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21o_1
X_185_ _057_ _048_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2_2
X_254_ u_uart.u_tx.clk_cnt\[13\] _108_ net10 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload2 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_EDGE_ROW_28_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ cpu_acc\[6\] _133_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand2_1
X_237_ _098_ _099_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nor2_1
Xhold14 u_uart.tx_data\[7\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 cpu_pc\[0\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 u_uart.u_tx.clk_cnt\[5\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_270_ cpu_pc\[1\] cpu_acc\[1\] _059_ _063_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__or4_1
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_399_ clknet_3_2__leaf_clk _016_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_322_ u_uart.tx_data\[2\] _158_ net8 net63 VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__a22o_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_184_ net30 _062_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nor2_1
X_253_ _108_ _109_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_2
X_305_ cpu_acc\[6\] _133_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_3_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_236_ net50 _096_ _083_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold26 u_uart.tx_data\[3\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold15 _032_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold37 u_uart.u_tx.clk_cnt\[10\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_219_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] u_uart.u_tx.clk_cnt\[2\]
+ net10 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a31o_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_398_ clknet_3_2__leaf_clk _015_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_321_ net25 _160_ _163_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__a21o_1
X_183_ u_cpu.state\[0\] _061_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_252_ net52 _107_ _083_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__o21ai_1
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__bufinv_16
X_304_ _141_ _145_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__and3_1
X_235_ u_uart.u_tx.clk_cnt\[5\] u_uart.u_tx.clk_cnt\[4\] u_uart.u_tx.clk_cnt\[6\]
+ _088_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__and4_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold16 u_uart.u_tx.shifter\[3\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 u_uart.tx_data\[2\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 u_uart.u_tx.clk_cnt\[13\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_218_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] u_uart.u_tx.clk_cnt\[2\]
+ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_397_ clknet_3_3__leaf_clk _014_ net13 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_320_ u_uart.tx_data\[1\] _158_ _159_ net21 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__a22o_1
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_251_ u_uart.u_tx.clk_cnt\[12\] _107_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__and2_1
X_182_ _059_ _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nor2_1
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/X sky130_fd_sc_hd__clkbuf_8
X_303_ _132_ _134_ _135_ _142_ _146_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__a2111o_1
X_234_ _096_ _097_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__nor2_1
Xhold17 _028_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 cpu_acc\[3\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 u_uart.tx_data\[1\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ net61 net48 _084_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__o21a_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_396_ clknet_3_3__leaf_clk _013_ net13 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ net10 _106_ _107_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nor3_1
X_181_ cpu_pc\[1\] cpu_pc\[0\] cpu_pc\[3\] cpu_pc\[2\] VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__or4b_1
X_379_ clknet_3_7__leaf_clk net29 net17 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/X sky130_fd_sc_hd__clkbuf_4
X_302_ cpu_acc\[5\] _116_ net7 _148_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a22o_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ net54 _094_ _083_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 u_uart.tx_data\[0\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 cpu_pc\[4\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_216_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] net10 VGND VGND VPWR VPWR
+ _084_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_17_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_395_ clknet_3_3__leaf_clk _012_ net13 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout10 _082_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
X_180_ cpu_pc\[5\] cpu_pc\[4\] cpu_pc\[7\] cpu_pc\[6\] VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or4_2
X_378_ clknet_3_7__leaf_clk net35 net16 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_301_ _146_ _147_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_232_ u_uart.u_tx.clk_cnt\[5\] u_uart.u_tx.clk_cnt\[4\] _088_ VGND VGND VPWR VPWR
+ _096_ sky130_fd_sc_hd__and3_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold19 u_uart.tx_data\[5\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_215_ net48 net10 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nor2_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_394_ clknet_3_2__leaf_clk _011_ net13 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout11 net14 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
X_377_ clknet_3_7__leaf_clk _027_ net16 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ _140_ _143_ _141_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__o21ai_1
X_231_ u_uart.u_tx.clk_cnt\[4\] _088_ _093_ _095_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o211a_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 rst_n VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_10_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_214_ u_uart.u_tx.state\[1\] u_uart.u_tx.state\[0\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__or2_2
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_393_ clknet_3_2__leaf_clk _010_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout12 net14 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
X_376_ clknet_3_7__leaf_clk _026_ net16 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_230_ _082_ _094_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__nor2_1
X_359_ clknet_3_1__leaf_clk u_cpu.pc_next\[0\] net11 VGND VGND VPWR VPWR cpu_pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ u_uart.u_tx.state\[1\] u_uart.u_tx.state\[0\] VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nor2_1
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_392_ clknet_3_2__leaf_clk _009_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout13 net14 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_375_ clknet_3_6__leaf_clk _025_ net16 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_358_ _054_ _062_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and2_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ _132_ _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nand2_1
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ net20 _080_ VGND VGND VPWR VPWR u_cpu.pc_next\[7\] sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_27_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_391_ clknet_3_2__leaf_clk _008_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout14 net1 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_374_ clknet_3_4__leaf_clk _024_ net15 VGND VGND VPWR VPWR cpu_acc\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_288_ _134_ _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nand2_1
X_357_ net32 cpu_acc\[7\] _000_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__mux2_1
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_211_ _080_ _081_ VGND VGND VPWR VPWR u_cpu.pc_next\[6\] sky130_fd_sc_hd__and2_1
X_409_ clknet_3_4__leaf_clk _041_ net15 VGND VGND VPWR VPWR u_uart.tx_data\[2\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ clknet_3_2__leaf_clk _001_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout15 net18 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_373_ clknet_3_4__leaf_clk _023_ net15 VGND VGND VPWR VPWR cpu_acc\[6\] sky130_fd_sc_hd__dfrtp_1
X_356_ net41 cpu_acc\[6\] _000_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__mux2_1
X_287_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__inv_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_408_ clknet_3_6__leaf_clk _040_ net16 VGND VGND VPWR VPWR u_uart.tx_data\[1\] sky130_fd_sc_hd__dfrtp_1
X_210_ cpu_pc\[6\] _078_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__or2_1
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_339_ _093_ _172_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__nor2_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout16 net18 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
X_372_ clknet_3_5__leaf_clk _022_ net15 VGND VGND VPWR VPWR cpu_acc\[5\] sky130_fd_sc_hd__dfrtp_2
X_355_ net37 cpu_acc\[5\] _000_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__mux2_1
X_286_ cpu_acc\[3\] _133_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__nor2_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_338_ u_uart.u_tx.bit_cnt\[1\] u_uart.u_tx.bit_cnt\[0\] u_uart.u_tx.bit_cnt\[2\]
+ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__nand3_1
X_407_ clknet_3_6__leaf_clk _039_ net16 VGND VGND VPWR VPWR u_uart.tx_data\[0\] sky130_fd_sc_hd__dfrtp_1
X_269_ cpu_pc\[1\] _064_ cpu_acc\[1\] VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ clknet_3_5__leaf_clk _021_ net15 VGND VGND VPWR VPWR cpu_acc\[4\] sky130_fd_sc_hd__dfrtp_2
Xfanout17 net18 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_354_ net40 cpu_acc\[4\] _000_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__mux2_1
X_285_ cpu_acc\[3\] _133_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__nand2_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_337_ u_uart.u_tx.bit_cnt\[1\] u_uart.u_tx.bit_cnt\[0\] _161_ u_uart.u_tx.bit_cnt\[2\]
+ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__a31o_1
X_406_ clknet_3_6__leaf_clk _000_ net13 VGND VGND VPWR VPWR u_uart.tx_start sky130_fd_sc_hd__dfrtp_1
X_199_ cpu_pc\[1\] cpu_pc\[0\] cpu_pc\[2\] VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__and3_1
X_268_ cpu_pc\[1\] _059_ _063_ cpu_acc\[1\] VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o31a_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout18 net1 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
X_370_ clknet_3_4__leaf_clk _020_ net15 VGND VGND VPWR VPWR cpu_acc\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_353_ net44 cpu_acc\[3\] _000_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__mux2_1
X_284_ _064_ _071_ _061_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__o21ba_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_336_ _169_ _170_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nor2_1
X_267_ cpu_acc\[0\] _116_ _118_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a21o_1
X_405_ clknet_3_0__leaf_clk _007_ net11 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_198_ _070_ _073_ VGND VGND VPWR VPWR u_cpu.pc_next\[1\] sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_319_ _162_ net36 net9 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_352_ net45 cpu_acc\[2\] _000_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__mux2_1
X_283_ _128_ _130_ _127_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o21ba_1
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_335_ u_uart.u_tx.bit_cnt\[1\] u_uart.u_tx.bit_cnt\[0\] net8 _158_ VGND VGND VPWR
+ VPWR _170_ sky130_fd_sc_hd__a31o_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_266_ u_cpu.state\[0\] _054_ _058_ _073_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__o221a_1
X_404_ clknet_3_0__leaf_clk _006_ net11 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_197_ _071_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_318_ u_uart.u_tx.shifter\[0\] u_uart.u_tx.shifter\[1\] net8 VGND VGND VPWR VPWR
+ _162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ u_uart.u_tx.clk_cnt\[11\] u_uart.u_tx.clk_cnt\[10\] _103_ VGND VGND VPWR VPWR
+ _107_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 u_uart.u_tx.clk_cnt\[15\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_420_ cpu_acc\[3\] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_282_ _124_ _131_ cpu_acc\[2\] _117_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__o2bb2a_1
X_351_ net46 cpu_acc\[1\] _000_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__mux2_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_334_ u_uart.u_tx.bit_cnt\[0\] _161_ net59 VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__a21oi_1
X_403_ clknet_3_0__leaf_clk _005_ net11 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__inv_2
X_196_ cpu_pc\[1\] _055_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nor2_1
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_317_ net9 net8 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__or2_1
X_179_ cpu_acc\[0\] VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__inv_2
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ u_uart.u_tx.clk_cnt\[10\] _103_ u_uart.u_tx.clk_cnt\[11\] VGND VGND VPWR VPWR
+ _106_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 cpu_pc\[7\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_350_ net36 cpu_acc\[0\] _000_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
X_281_ _129_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__xor2_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_333_ net8 _160_ u_uart.u_tx.bit_cnt\[0\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__mux2_1
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_264_ _065_ _067_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or2_4
X_402_ clknet_3_2__leaf_clk _004_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_195_ cpu_pc\[1\] _055_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_316_ net9 net8 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_26_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ net55 _103_ _105_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o21a_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_178_ u_uart.tx_busy VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3 u_uart.u_tx.shifter\[2\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_280_ _121_ _122_ _119_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_332_ net32 net9 _160_ u_uart.u_tx.shifter\[7\] VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a22o_1
X_263_ net24 _115_ _114_ VGND VGND VPWR VPWR u_uart.u_tx.tx_next sky130_fd_sc_hd__o21a_1
X_401_ clknet_3_2__leaf_clk _003_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_194_ net43 _070_ VGND VGND VPWR VPWR u_cpu.pc_next\[0\] sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_315_ _093_ _115_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__nor2_1
X_177_ u_uart.u_tx.state\[0\] VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__inv_2
X_246_ u_uart.u_tx.clk_cnt\[10\] _103_ net10 VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ u_uart.u_tx.clk_cnt\[4\] _088_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__and2_1
Xhold4 u_uart.u_tx.shifter\[5\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ net26 _160_ _168_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21o_1
X_262_ u_uart.u_tx.state\[1\] _056_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__nand2_1
X_193_ _065_ _066_ _068_ _069_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or4_1
X_400_ clknet_3_2__leaf_clk _002_ net12 VGND VGND VPWR VPWR u_uart.u_tx.clk_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_314_ u_uart.tx_start _057_ net10 VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__and3_1
X_245_ _103_ _104_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nor2_1
X_176_ cpu_pc\[0\] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
XFILLER_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_228_ _089_ _090_ _091_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__or4_4
XFILLER_17_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 _030_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ u_uart.tx_data\[6\] net9 net8 u_uart.u_tx.shifter\[7\] VGND VGND VPWR VPWR
+ _168_ sky130_fd_sc_hd__a22o_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_261_ u_uart.u_tx.state\[1\] _056_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__or2_1
X_192_ cpu_acc\[1\] cpu_acc\[0\] cpu_acc\[2\] cpu_acc\[3\] VGND VGND VPWR VPWR _069_
+ sky130_fd_sc_hd__or4_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_313_ net38 _116_ net7 _157_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a22o_1
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_175_ u_cpu.state\[1\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__inv_2
X_244_ net53 _102_ _083_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ u_uart.u_tx.clk_cnt\[5\] u_uart.u_tx.clk_cnt\[4\] u_uart.u_tx.clk_cnt\[7\]
+ u_uart.u_tx.clk_cnt\[6\] VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__or4_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 u_uart.u_tx.shifter\[0\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_260_ net19 _112_ _113_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
X_389_ clknet_3_6__leaf_clk _038_ net16 VGND VGND VPWR VPWR u_uart.u_tx.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_191_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__inv_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_312_ _155_ _156_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_243_ u_uart.u_tx.clk_cnt\[7\] u_uart.u_tx.clk_cnt\[9\] u_uart.u_tx.clk_cnt\[8\]
+ _098_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_226_ u_uart.u_tx.clk_cnt\[9\] u_uart.u_tx.clk_cnt\[8\] u_uart.u_tx.clk_cnt\[11\]
+ u_uart.u_tx.clk_cnt\[10\] VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__or4_1
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 u_uart.u_tx.shifter\[1\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
X_209_ cpu_pc\[6\] _078_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand2_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ cpu_pc\[1\] cpu_pc\[0\] VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__and2_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_388_ clknet_3_3__leaf_clk _037_ net12 VGND VGND VPWR VPWR u_uart.u_tx.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ cpu_acc\[7\] _133_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__xor2_1
XFILLER_14_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_242_ net10 _101_ _102_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_21_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ u_uart.u_tx.clk_cnt\[13\] u_uart.u_tx.clk_cnt\[12\] u_uart.u_tx.clk_cnt\[15\]
+ u_uart.u_tx.clk_cnt\[14\] VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__or4_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 u_uart.u_tx.shifter\[6\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_208_ _078_ _079_ VGND VGND VPWR VPWR u_cpu.pc_next\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_387_ clknet_3_6__leaf_clk _036_ net16 VGND VGND VPWR VPWR u_uart.tx_busy sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _141_ _145_ _149_ _152_ _151_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__a41o_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ u_uart.u_tx.clk_cnt\[7\] u_uart.u_tx.clk_cnt\[8\] _098_ VGND VGND VPWR VPWR
+ _102_ sky130_fd_sc_hd__and3_1
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_224_ _083_ _087_ _089_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and3_1
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold9 _031_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_207_ net62 _076_ net42 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire7 _126_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_386_ clknet_3_7__leaf_clk u_uart.u_tx.tx_next net16 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfstp_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_240_ u_uart.u_tx.clk_cnt\[7\] _098_ u_uart.u_tx.clk_cnt\[8\] VGND VGND VPWR VPWR
+ _101_ sky130_fd_sc_hd__a21oi_1
X_369_ clknet_3_4__leaf_clk _019_ net15 VGND VGND VPWR VPWR cpu_acc\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_223_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] u_uart.u_tx.clk_cnt\[3\]
+ u_uart.u_tx.clk_cnt\[2\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand4_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_206_ cpu_pc\[5\] cpu_pc\[4\] _076_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__and3_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_385_ clknet_3_7__leaf_clk _035_ net17 VGND VGND VPWR VPWR u_uart.u_tx.bit_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_299_ cpu_acc\[5\] _133_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__xnor2_1
X_368_ clknet_3_1__leaf_clk _018_ net14 VGND VGND VPWR VPWR cpu_acc\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_222_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] u_uart.u_tx.clk_cnt\[3\]
+ u_uart.u_tx.clk_cnt\[2\] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__and4_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ net47 _076_ VGND VGND VPWR VPWR u_cpu.pc_next\[4\] sky130_fd_sc_hd__xor2_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_384_ clknet_3_7__leaf_clk _034_ net17 VGND VGND VPWR VPWR u_uart.u_tx.bit_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput2 net2 VGND VGND VPWR VPWR gpio[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ cpu_acc\[5\] _133_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__nand2_1
X_367_ clknet_3_4__leaf_clk _017_ net15 VGND VGND VPWR VPWR cpu_acc\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ u_uart.u_tx.clk_cnt\[1\] u_uart.u_tx.clk_cnt\[0\] u_uart.u_tx.clk_cnt\[2\]
+ u_uart.u_tx.clk_cnt\[3\] VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__a31o_1
X_419_ cpu_acc\[2\] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_204_ _076_ _077_ VGND VGND VPWR VPWR u_cpu.pc_next\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_383_ clknet_3_7__leaf_clk _033_ net17 VGND VGND VPWR VPWR u_uart.u_tx.bit_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput3 net3 VGND VGND VPWR VPWR gpio[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_297_ cpu_acc\[4\] _116_ net7 _144_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a22o_1
X_366_ clknet_3_0__leaf_clk u_cpu.pc_next\[7\] net11 VGND VGND VPWR VPWR cpu_pc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_220_ _085_ _086_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__nor2_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ _093_ _114_ _053_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__o21ai_1
X_418_ cpu_acc\[1\] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_203_ net49 _074_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nor2_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ clknet_3_6__leaf_clk net33 net16 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput4 net4 VGND VGND VPWR VPWR gpio[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ _142_ _143_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__xor2_1
XFILLER_13_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_365_ clknet_3_0__leaf_clk u_cpu.pc_next\[6\] net11 VGND VGND VPWR VPWR cpu_pc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ net51 _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_279_ _127_ _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nor2_1
X_417_ cpu_acc\[0\] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_29_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_202_ cpu_pc\[3\] _074_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR gpio[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_381_ clknet_3_7__leaf_clk net27 net17 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_295_ _132_ _134_ _135_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__a21o_1
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_364_ clknet_3_0__leaf_clk u_cpu.pc_next\[5\] net11 VGND VGND VPWR VPWR cpu_pc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_347_ _115_ _173_ _051_ _052_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__o211a_1
X_278_ _055_ cpu_acc\[2\] _064_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nor3_1
X_416_ clknet_3_6__leaf_clk net31 net13 VGND VGND VPWR VPWR u_cpu.state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_201_ _074_ _075_ VGND VGND VPWR VPWR u_cpu.pc_next\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 cpu_pc\[2\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_380_ clknet_3_7__leaf_clk net23 net17 VGND VGND VPWR VPWR u_uart.u_tx.shifter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput6 net6 VGND VGND VPWR VPWR uart_tx sky130_fd_sc_hd__buf_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

